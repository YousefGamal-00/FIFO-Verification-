package shared_pkg_0;

bit test_finished; 
int error_count; 
int correct_count;

endpackage